module virp
