module vrpc
