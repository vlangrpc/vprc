module vrpc

pub enum ErrorCode {
	ok    = 0
	error = 1
}
